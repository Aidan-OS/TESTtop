Club|false|0|0|A generic club.|Light|2|0.1|1d4*Bludgeoning|