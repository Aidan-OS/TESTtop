Javelin|false|0|0|A generic javelin.|Thrown (range 30/120)|2|0.5|1d6*Piercing|