Dagger|false|0|0|A generic dagger.|Finesse, Light, Thrown (range 20/60)|1|2|1d4*Piercing|